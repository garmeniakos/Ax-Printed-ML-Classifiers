//weights: [[[40, -34, 40, 20, 8, -4, 76, 32, 28, -34, -42, 8, -60, -24, 28, 28, -32, -48, -48, 68, -15], [-12, -8, -15, -16, -4, 28, 16, 32, 12, 48, 8, 28, 16, 4, -24, 1, 2, 20, -40, 9, 0], [28, -56, 36, -34, 0, 16, 48, 48, -4, 18, -24, -24, -4, 18, 16, -24, -32, -7, 16, 12, 8]], [[44, 60, 48]]]
//intercepts: [[370, 187, -222], [37311]]
//act size: [4, 13, 21]
//pred num: 1
module top (inp, out);
input [83:0] inp;
output [21:0] out;

// layer: 0 - neuron: 0
    wire signed [11:0] n_0_0_po_0;
    //weight 40: 8'sb00101000
    assign n_0_0_po_0 = $signed({1'b0, inp[3:0]}) * 8'sb00101000;

    wire signed [11:0] n_0_0_po_1;
    //weight -34: 8'sb11011110
    assign n_0_0_po_1 = $signed({1'b0, inp[7:4]}) * 8'sb11011110;

    wire signed [11:0] n_0_0_po_2;
    //weight 40: 8'sb00101000
    assign n_0_0_po_2 = $signed({1'b0, inp[11:8]}) * 8'sb00101000;

    wire signed [11:0] n_0_0_po_3;
    //weight 20: 8'sb00010100
    assign n_0_0_po_3 = $signed({1'b0, inp[15:12]}) * 8'sb00010100;

    wire signed [11:0] n_0_0_po_4;
    //weight 8: 8'sb00001000
    assign n_0_0_po_4 = $signed({1'b0, inp[19:16]}) * 8'sb00001000;

    wire signed [11:0] n_0_0_po_5;
    //weight -4: 8'sb11111100
    assign n_0_0_po_5 = $signed({1'b0, inp[23:20]}) * 8'sb11111100;

    wire signed [11:0] n_0_0_po_6;
    //weight 76: 8'sb01001100
    assign n_0_0_po_6 = $signed({1'b0, inp[27:24]}) * 8'sb01001100;

    wire signed [11:0] n_0_0_po_7;
    //weight 32: 8'sb00100000
    assign n_0_0_po_7 = $signed({1'b0, inp[31:28]}) * 8'sb00100000;

    wire signed [11:0] n_0_0_po_8;
    //weight 28: 8'sb00011100
    assign n_0_0_po_8 = $signed({1'b0, inp[35:32]}) * 8'sb00011100;

    wire signed [11:0] n_0_0_po_9;
    //weight -34: 8'sb11011110
    assign n_0_0_po_9 = $signed({1'b0, inp[39:36]}) * 8'sb11011110;

    wire signed [11:0] n_0_0_po_10;
    //weight -42: 8'sb11010110
    assign n_0_0_po_10 = $signed({1'b0, inp[43:40]}) * 8'sb11010110;

    wire signed [11:0] n_0_0_po_11;
    //weight 8: 8'sb00001000
    assign n_0_0_po_11 = $signed({1'b0, inp[47:44]}) * 8'sb00001000;

    wire signed [11:0] n_0_0_po_12;
    //weight -60: 8'sb11000100
    assign n_0_0_po_12 = $signed({1'b0, inp[51:48]}) * 8'sb11000100;

    wire signed [11:0] n_0_0_po_13;
    //weight -24: 8'sb11101000
    assign n_0_0_po_13 = $signed({1'b0, inp[55:52]}) * 8'sb11101000;

    wire signed [11:0] n_0_0_po_14;
    //weight 28: 8'sb00011100
    assign n_0_0_po_14 = $signed({1'b0, inp[59:56]}) * 8'sb00011100;

    wire signed [11:0] n_0_0_po_15;
    //weight 28: 8'sb00011100
    assign n_0_0_po_15 = $signed({1'b0, inp[63:60]}) * 8'sb00011100;

    wire signed [11:0] n_0_0_po_16;
    //weight -32: 8'sb11100000
    assign n_0_0_po_16 = $signed({1'b0, inp[67:64]}) * 8'sb11100000;

    wire signed [11:0] n_0_0_po_17;
    //weight -48: 8'sb11010000
    assign n_0_0_po_17 = $signed({1'b0, inp[71:68]}) * 8'sb11010000;

    wire signed [11:0] n_0_0_po_18;
    //weight -48: 8'sb11010000
    assign n_0_0_po_18 = $signed({1'b0, inp[75:72]}) * 8'sb11010000;

    wire signed [11:0] n_0_0_po_19;
    //weight 68: 8'sb01000100
    assign n_0_0_po_19 = $signed({1'b0, inp[79:76]}) * 8'sb01000100;

    wire signed [11:0] n_0_0_po_20;
    //weight -15: 8'sb11110001
    assign n_0_0_po_20 = $signed({1'b0, inp[83:80]}) * 8'sb11110001;

    wire signed [13:0] n_0_0_sum;
    assign n_0_0_sum = 370 + n_0_0_po_0 + n_0_0_po_1 + n_0_0_po_2 + n_0_0_po_3 + n_0_0_po_4 + n_0_0_po_5 + n_0_0_po_6 + n_0_0_po_7 + n_0_0_po_8 + n_0_0_po_9 + n_0_0_po_10 + n_0_0_po_11 + n_0_0_po_12 + n_0_0_po_13 + n_0_0_po_14 + n_0_0_po_15 + n_0_0_po_16 + n_0_0_po_17 + n_0_0_po_18 + n_0_0_po_19 + n_0_0_po_20;
    //relu
    wire [12:0] n_0_0;
    assign n_0_0 = (n_0_0_sum<0) ? $unsigned({13{1'b0}}) : $unsigned(n_0_0_sum[12:0]);

// layer: 0 - neuron: 1
    wire signed [11:0] n_0_1_po_0;
    //weight -12: 8'sb11110100
    assign n_0_1_po_0 = $signed({1'b0, inp[3:0]}) * 8'sb11110100;

    wire signed [11:0] n_0_1_po_1;
    //weight -8: 8'sb11111000
    assign n_0_1_po_1 = $signed({1'b0, inp[7:4]}) * 8'sb11111000;

    wire signed [11:0] n_0_1_po_2;
    //weight -15: 8'sb11110001
    assign n_0_1_po_2 = $signed({1'b0, inp[11:8]}) * 8'sb11110001;

    wire signed [11:0] n_0_1_po_3;
    //weight -16: 8'sb11110000
    assign n_0_1_po_3 = $signed({1'b0, inp[15:12]}) * 8'sb11110000;

    wire signed [11:0] n_0_1_po_4;
    //weight -4: 8'sb11111100
    assign n_0_1_po_4 = $signed({1'b0, inp[19:16]}) * 8'sb11111100;

    wire signed [11:0] n_0_1_po_5;
    //weight 28: 8'sb00011100
    assign n_0_1_po_5 = $signed({1'b0, inp[23:20]}) * 8'sb00011100;

    wire signed [11:0] n_0_1_po_6;
    //weight 16: 8'sb00010000
    assign n_0_1_po_6 = $signed({1'b0, inp[27:24]}) * 8'sb00010000;

    wire signed [11:0] n_0_1_po_7;
    //weight 32: 8'sb00100000
    assign n_0_1_po_7 = $signed({1'b0, inp[31:28]}) * 8'sb00100000;

    wire signed [11:0] n_0_1_po_8;
    //weight 12: 8'sb00001100
    assign n_0_1_po_8 = $signed({1'b0, inp[35:32]}) * 8'sb00001100;

    wire signed [11:0] n_0_1_po_9;
    //weight 48: 8'sb00110000
    assign n_0_1_po_9 = $signed({1'b0, inp[39:36]}) * 8'sb00110000;

    wire signed [11:0] n_0_1_po_10;
    //weight 8: 8'sb00001000
    assign n_0_1_po_10 = $signed({1'b0, inp[43:40]}) * 8'sb00001000;

    wire signed [11:0] n_0_1_po_11;
    //weight 28: 8'sb00011100
    assign n_0_1_po_11 = $signed({1'b0, inp[47:44]}) * 8'sb00011100;

    wire signed [11:0] n_0_1_po_12;
    //weight 16: 8'sb00010000
    assign n_0_1_po_12 = $signed({1'b0, inp[51:48]}) * 8'sb00010000;

    wire signed [11:0] n_0_1_po_13;
    //weight 4: 8'sb00000100
    assign n_0_1_po_13 = $signed({1'b0, inp[55:52]}) * 8'sb00000100;

    wire signed [11:0] n_0_1_po_14;
    //weight -24: 8'sb11101000
    assign n_0_1_po_14 = $signed({1'b0, inp[59:56]}) * 8'sb11101000;

    wire signed [11:0] n_0_1_po_15;
    //weight 1: 8'sb00000001
    assign n_0_1_po_15 = $signed({1'b0, inp[63:60]}) * 8'sb00000001;

    wire signed [11:0] n_0_1_po_16;
    //weight 2: 8'sb00000010
    assign n_0_1_po_16 = $signed({1'b0, inp[67:64]}) * 8'sb00000010;

    wire signed [11:0] n_0_1_po_17;
    //weight 20: 8'sb00010100
    assign n_0_1_po_17 = $signed({1'b0, inp[71:68]}) * 8'sb00010100;

    wire signed [11:0] n_0_1_po_18;
    //weight -40: 8'sb11011000
    assign n_0_1_po_18 = $signed({1'b0, inp[75:72]}) * 8'sb11011000;

    wire signed [11:0] n_0_1_po_19;
    //weight 9: 8'sb00001001
    assign n_0_1_po_19 = $signed({1'b0, inp[79:76]}) * 8'sb00001001;

    wire signed [11:0] n_0_1_po_20;
    //weight 0: 8'sb00000000
    assign n_0_1_po_20 = $signed({1'b0, inp[83:80]}) * 8'sb00000000;

    wire signed [13:0] n_0_1_sum;
    assign n_0_1_sum = 187 + n_0_1_po_0 + n_0_1_po_1 + n_0_1_po_2 + n_0_1_po_3 + n_0_1_po_4 + n_0_1_po_5 + n_0_1_po_6 + n_0_1_po_7 + n_0_1_po_8 + n_0_1_po_9 + n_0_1_po_10 + n_0_1_po_11 + n_0_1_po_12 + n_0_1_po_13 + n_0_1_po_14 + n_0_1_po_15 + n_0_1_po_16 + n_0_1_po_17 + n_0_1_po_18 + n_0_1_po_19 + n_0_1_po_20;
    //relu
    wire [12:0] n_0_1;
    assign n_0_1 = (n_0_1_sum<0) ? $unsigned({13{1'b0}}) : $unsigned(n_0_1_sum[12:0]);

// layer: 0 - neuron: 2
    wire signed [11:0] n_0_2_po_0;
    //weight 28: 8'sb00011100
    assign n_0_2_po_0 = $signed({1'b0, inp[3:0]}) * 8'sb00011100;

    wire signed [11:0] n_0_2_po_1;
    //weight -56: 8'sb11001000
    assign n_0_2_po_1 = $signed({1'b0, inp[7:4]}) * 8'sb11001000;

    wire signed [11:0] n_0_2_po_2;
    //weight 36: 8'sb00100100
    assign n_0_2_po_2 = $signed({1'b0, inp[11:8]}) * 8'sb00100100;

    wire signed [11:0] n_0_2_po_3;
    //weight -34: 8'sb11011110
    assign n_0_2_po_3 = $signed({1'b0, inp[15:12]}) * 8'sb11011110;

    wire signed [11:0] n_0_2_po_4;
    //weight 0: 8'sb00000000
    assign n_0_2_po_4 = $signed({1'b0, inp[19:16]}) * 8'sb00000000;

    wire signed [11:0] n_0_2_po_5;
    //weight 16: 8'sb00010000
    assign n_0_2_po_5 = $signed({1'b0, inp[23:20]}) * 8'sb00010000;

    wire signed [11:0] n_0_2_po_6;
    //weight 48: 8'sb00110000
    assign n_0_2_po_6 = $signed({1'b0, inp[27:24]}) * 8'sb00110000;

    wire signed [11:0] n_0_2_po_7;
    //weight 48: 8'sb00110000
    assign n_0_2_po_7 = $signed({1'b0, inp[31:28]}) * 8'sb00110000;

    wire signed [11:0] n_0_2_po_8;
    //weight -4: 8'sb11111100
    assign n_0_2_po_8 = $signed({1'b0, inp[35:32]}) * 8'sb11111100;

    wire signed [11:0] n_0_2_po_9;
    //weight 18: 8'sb00010010
    assign n_0_2_po_9 = $signed({1'b0, inp[39:36]}) * 8'sb00010010;

    wire signed [11:0] n_0_2_po_10;
    //weight -24: 8'sb11101000
    assign n_0_2_po_10 = $signed({1'b0, inp[43:40]}) * 8'sb11101000;

    wire signed [11:0] n_0_2_po_11;
    //weight -24: 8'sb11101000
    assign n_0_2_po_11 = $signed({1'b0, inp[47:44]}) * 8'sb11101000;

    wire signed [11:0] n_0_2_po_12;
    //weight -4: 8'sb11111100
    assign n_0_2_po_12 = $signed({1'b0, inp[51:48]}) * 8'sb11111100;

    wire signed [11:0] n_0_2_po_13;
    //weight 18: 8'sb00010010
    assign n_0_2_po_13 = $signed({1'b0, inp[55:52]}) * 8'sb00010010;

    wire signed [11:0] n_0_2_po_14;
    //weight 16: 8'sb00010000
    assign n_0_2_po_14 = $signed({1'b0, inp[59:56]}) * 8'sb00010000;

    wire signed [11:0] n_0_2_po_15;
    //weight -24: 8'sb11101000
    assign n_0_2_po_15 = $signed({1'b0, inp[63:60]}) * 8'sb11101000;

    wire signed [11:0] n_0_2_po_16;
    //weight -32: 8'sb11100000
    assign n_0_2_po_16 = $signed({1'b0, inp[67:64]}) * 8'sb11100000;

    wire signed [11:0] n_0_2_po_17;
    //weight -7: 8'sb11111001
    assign n_0_2_po_17 = $signed({1'b0, inp[71:68]}) * 8'sb11111001;

    wire signed [11:0] n_0_2_po_18;
    //weight 16: 8'sb00010000
    assign n_0_2_po_18 = $signed({1'b0, inp[75:72]}) * 8'sb00010000;

    wire signed [11:0] n_0_2_po_19;
    //weight 12: 8'sb00001100
    assign n_0_2_po_19 = $signed({1'b0, inp[79:76]}) * 8'sb00001100;

    wire signed [11:0] n_0_2_po_20;
    //weight 8: 8'sb00001000
    assign n_0_2_po_20 = $signed({1'b0, inp[83:80]}) * 8'sb00001000;

    wire signed [13:0] n_0_2_sum;
    assign n_0_2_sum = -222 + n_0_2_po_0 + n_0_2_po_1 + n_0_2_po_2 + n_0_2_po_3 + n_0_2_po_4 + n_0_2_po_5 + n_0_2_po_6 + n_0_2_po_7 + n_0_2_po_8 + n_0_2_po_9 + n_0_2_po_10 + n_0_2_po_11 + n_0_2_po_12 + n_0_2_po_13 + n_0_2_po_14 + n_0_2_po_15 + n_0_2_po_16 + n_0_2_po_17 + n_0_2_po_18 + n_0_2_po_19 + n_0_2_po_20;
    //relu
    wire [12:0] n_0_2;
    assign n_0_2 = (n_0_2_sum<0) ? $unsigned({13{1'b0}}) : $unsigned(n_0_2_sum[12:0]);

// layer: 1 - neuron: 0
    wire signed [20:0] n_1_0_po_0;
    //weight 44: 8'sb00101100
    assign n_1_0_po_0 = $signed({1'b0, n_0_0}) * 8'sb00101100;

    wire signed [20:0] n_1_0_po_1;
    //weight 60: 8'sb00111100
    assign n_1_0_po_1 = $signed({1'b0, n_0_1}) * 8'sb00111100;

    wire signed [20:0] n_1_0_po_2;
    //weight 48: 8'sb00110000
    assign n_1_0_po_2 = $signed({1'b0, n_0_2}) * 8'sb00110000;

    wire signed [21:0] n_1_0_sum;
    assign n_1_0_sum = 37311 + n_1_0_po_0 + n_1_0_po_1 + n_1_0_po_2;
    //relu
    wire [20:0] n_1_0;
    assign n_1_0 = (n_1_0_sum<0) ? $unsigned({21{1'b0}}) : $unsigned(n_1_0_sum[20:0]);

    assign out = {n_1_0};

endmodule
